//inside TB module
import "DPI-C" context function void function_name();
// use imported function in SystemVerilog
// export "DPI-C" context task sv_function_name();
// use exported function in C
